LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY driver7Segmentos IS
 PORT( codigoCaracter : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
 bitsCaracter : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END driver7Segmentos;
ARCHITECTURE Structure OF driver7Segmentos IS
BEGIN
 .
. -- Aquí debéis poner vuestro código que implemente el driver
.
END Structure;